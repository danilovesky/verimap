module empty (i, z);
  input i;
  output z;
  BU1 inst_z (.A(i), .Q(z));
endmodule

module spinv1 (i, z);
  input i;
  output z;
  BU1 inst_z (.A(i), .Q(z));
endmodule

module spinv2 (i, z);
  input i;
  output z;
  BU1 inst_z (.A(i), .Q(z));
endmodule

module spinv3 (i, z);
  input i;
  output z;
  BU1 inst_z (.A(i), .Q(z));
endmodule

module spinv4 (i, z);
  input i;
  output z;
  BU1 inst_z (.A(i), .Q(z));
endmodule

module spinv8 (i, z);
  input i;
  output z;
  BU1 inst_z (.A(i), .Q(z));
endmodule
